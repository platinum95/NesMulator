`timescale 1ns / 1ps

package Common;

typedef struct {
    shortint PC;
    byte A, X, Y, S;
    byte P;
} CPUState;

endpackage
